LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use std.textio.all;
use work.txt_util.all;

entity execute_tb is
end execute_tb;
